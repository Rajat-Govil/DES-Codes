module IP_inv(
    input [1:64] round_in,
    output [1:64] ciphertext
    );
assign ciphertext[1] = round_in[40];
assign ciphertext[2] = round_in[8];
assign ciphertext[3] = round_in[48];
assign ciphertext[4] = round_in[16];
assign ciphertext[5] = round_in[56];
assign ciphertext[6] = round_in[24];
assign ciphertext[7] = round_in[64];
assign ciphertext[8] = round_in[32];
assign ciphertext[9] = round_in[39];
assign ciphertext[10] = round_in[7];
assign ciphertext[11] = round_in[47];
assign ciphertext[12] = round_in[15];
assign ciphertext[13] = round_in[55];
assign ciphertext[14] = round_in[23];
assign ciphertext[15] = round_in[63];
assign ciphertext[16] = round_in[31];
assign ciphertext[17] = round_in[38];
assign ciphertext[18] = round_in[6];
assign ciphertext[19] = round_in[46];
assign ciphertext[20] = round_in[14];
assign ciphertext[21] = round_in[54];
assign ciphertext[22] = round_in[22];
assign ciphertext[23] = round_in[62];
assign ciphertext[24] = round_in[30];
assign ciphertext[25] = round_in[37];
assign ciphertext[26] = round_in[5];
assign ciphertext[27] = round_in[45];
assign ciphertext[28] = round_in[13];
assign ciphertext[29] = round_in[53];
assign ciphertext[30] = round_in[21];
assign ciphertext[31] = round_in[61];
assign ciphertext[32] = round_in[29];
assign ciphertext[33] = round_in[36];
assign ciphertext[34] = round_in[4];
assign ciphertext[35] = round_in[44];
assign ciphertext[36] = round_in[12];
assign ciphertext[37] = round_in[52];
assign ciphertext[38] = round_in[20];
assign ciphertext[39] = round_in[60];
assign ciphertext[40] = round_in[28];
assign ciphertext[41] = round_in[35];
assign ciphertext[42] = round_in[3];
assign ciphertext[43] = round_in[43];
assign ciphertext[44] = round_in[11];
assign ciphertext[45] = round_in[51];
assign ciphertext[46] = round_in[19];
assign ciphertext[47] = round_in[59];
assign ciphertext[48] = round_in[27];
assign ciphertext[49] = round_in[34];
assign ciphertext[50] = round_in[2];
assign ciphertext[51] = round_in[42];
assign ciphertext[52] = round_in[10];
assign ciphertext[53] = round_in[50];
assign ciphertext[54] = round_in[18];
assign ciphertext[55] = round_in[58];
assign ciphertext[56] = round_in[26];
assign ciphertext[57] = round_in[33];
assign ciphertext[58] = round_in[1];
assign ciphertext[59] = round_in[41];
assign ciphertext[60] = round_in[9];
assign ciphertext[61] = round_in[49];
assign ciphertext[62] = round_in[17];
assign ciphertext[63] = round_in[57];
assign ciphertext[64] = round_in[25];
endmodule
